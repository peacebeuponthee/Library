* AD795 SPICE Macro-model        
* Description: Amplifier 
* Generic Desc: 8/30V, JFET, OP, Low Pwr, Low Noise, 1X
* Developed by: JOM / ADSC
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (11/1994)
* Copyright 1990, 2012 by Analog Devices.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*
* Parameters modeled include:
*
* END Notes
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD795    1 2 99 50 30
*
* INPUT STAGE & POLE AT 40 MHZ
*
R3   5  50    .719
R4   6  50    .719
CIN  1   2    2E-12
C2   5   6    1.383E-9
I1   99  4    100E-3
IOS  1   2    0.1E-12
EOS  65  1    POLY(1)  17 24  50E-6  1
J1   5   2    4   JX
J2   6   7    4   JX
EN   7  65    43  0  1
GN1  0   1    47  0  1E-6
GN2  0   2    61  0  1E-6
GB1  2  50    POLY(3) 4,2 5,2 50,2 0 1E-12 1E-12 1E-12
GB2  7  50    POLY(3) 4,7 6,7 50,7 0 1E-12 1E-12 1E-12
*
EREF 98  0    24  0   1
*
* VOLTAGE NOISE GENERATOR
*
VN1  41  0    DC 2
RS1  41 42    8E3
RS2  42 43    1.2E9
CS1  42 43    398E-11
RS3  43 44    1.2E9
CS2  43 44    398E-11
RS4  44 45    8E3
VN2  0  45    DC 2
*
* CURRENT NOISE GENERATOR
*
VN3  46  0    DC 2
RN5  46 47    41.5
RN6  47 48    41.5
VN4  0  48    DC 2
*
* CURRENT NOISE GENERATOR
*
VN5  60  0    DC 2
RN7  60 61    41.5
RN8  61 62    41.5
VN6  0  62    DC 2
*  
* SECOND STAGE & POLE AT 2.213 HZ
*
R5   9  98    719203
C3   9  98    1.00E-7
G1   98  9    5  6  1.39
V2   99  8    3.025
V3   10 50    3.025
D1   9   8    DX
D2   10  9    DX
*
* NEGATIVE ZERO AT 15 MHZ
*
R6   11 12     1E6
R7   12 98     1
E2   11 98     9  24  1E6
VX1  84  0    
EX1  83  0     11 12  1
FX1  11 12     VX1  -1
CX1  83 84     10.6E-15
*
* POLE AT 20 MHZ
*
R8   13 98     1E3
C5   13 98     7.96E-12
G2   98 13     12 24  1E-3
*
* POLE AT 20 MHZ
*
R9   14 98     1E3
C6   14 98     7.96E-12
G3   98 14     13 24  1E-3
*
* POLE AT 20 MHZ
*
R10  15 98     1E3
C7   15 98     7.96E-12
G4   98 15     14 24  1E-3
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 300 HZ
*
R11  16 17     1E6
C8   16 17     5.3E-10
R12  17 98     1
E3   16 98     POLY(2) 1  98  2  98  0  1.585  1.585
*
* POLE AT 20 MHZ
*
R13  18 98     1E3
C9   18 98     7.96E-12
G5   98 18     15 24  1E-3
*
* OUTPUT STAGE
*
R14  24 99     2000E3
R15  24 50     2000E3
FSY  99 50     POLY(2) V7 V8 -98.7E-3 1 1
R16  29 99     360
R17  29 50     360
L1   29 30     1E-8
G8   29 99     99 18  2.78E-3
G9   50 29     18 50  2.78E-3
V4   25 29     2.0
V5   29 26     2.0
D3   18 25     DX
D4   26 18     DX
F1   29  0     V4  1
F2   0  29     V5  1
G6   98 70     29 18 2.78E-3
D5   70 71     DX
D6   72 70     DX
V7   71 98     DC 0
V8   98 72     DC 0
*
* MODELS USED
*
.MODEL JX PJF(BETA=9.67  VTO=-2.000  IS=0.50E-12 RD=0.1
+ RS=0.1 CGD=1E-15 CGS=1E-15)
.MODEL DX   D(IS=1E-15 RS=10 CJO=1E-15)
.ENDS AD795


